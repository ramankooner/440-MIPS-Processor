`timescale 1ns / 1ps
/**********************************************************
*
*Author:   Raman Kooner, James Gojit
*Email:    ramankooner9@gmail.com, jamesjrgojit@gmail.com
*Filename: barrel_shifter.v
*Date:     November 20th, 2018
*Version:  1.3
*
*Notes: 
*
* The barrel shifter is used to shift a value by a certain 
* amount of bits. This allows us to use the shift amount
* field in our R-Type instructions. The barrel shifter is a
* case statement that looks for the shift type and will
* do a shift based on the amount of bits its being shifted.
*
***********************************************************/
module barrel_shifter(in, shift_type, shamt, out);

	// Inputs
	input  [31:0] in;
	input   [1:0] shift_type;
	input   [4:0] shamt;

	// Outupts and Registers
	output [31:0] out;
	reg    [31:0] out;

	always@(*) begin
		case({shift_type, shamt})
		
			//*******************************
			//************* KEY *************
			//*******************************
			
			//*******************************
			// SLL(I) - 00
			// SRL(I) - 01
			// SRA(I) - 10
			//*******************************
			
			// Shift Left Logical
			7'b00_00000: out = in[31:0];
			7'b00_00001: out = {in[30:0],1'b0 };
			7'b00_00010: out = {in[29:0],2'b0 };
			7'b00_00011: out = {in[28:0],3'b0 };
			7'b00_00100: out = {in[27:0],4'b0 };
			7'b00_00101: out = {in[26:0],5'b0 };
			7'b00_00110: out = {in[25:0],6'b0 };
			7'b00_00111: out = {in[24:0],7'b0 };
			7'b00_01000: out = {in[23:0],8'b0 };
			7'b00_01001: out = {in[22:0],9'b0 };
			7'b00_01010: out = {in[21:0],10'b0};
			7'b00_01011: out = {in[20:0],11'b0};
			7'b00_01100: out = {in[19:0],12'b0};
			7'b00_01101: out = {in[18:0],13'b0};
			7'b00_01110: out = {in[17:0],14'b0};
			7'b00_01111: out = {in[16:0],15'b0};
			7'b00_10000: out = {in[15:0],16'b0};
			7'b00_10001: out = {in[14:0],17'b0};
			7'b00_10010: out = {in[13:0],18'b0};
			7'b00_10011: out = {in[12:0],19'b0};
			7'b00_10100: out = {in[11:0],20'b0};
			7'b00_10101: out = {in[10:0],21'b0};
			7'b00_10110: out = { in[9:0],22'b0};
			7'b00_10111: out = { in[8:0],23'b0};
			7'b00_11000: out = { in[7:0],24'b0};
			7'b00_11001: out = { in[6:0],25'b0};
			7'b00_11010: out = { in[5:0],26'b0};
			7'b00_11011: out = { in[4:0],27'b0};
			7'b00_11100: out = { in[3:0],28'b0};
			7'b00_11101: out = { in[2:0],29'b0};
			7'b00_11110: out = { in[1:0],30'b0};
			7'b00_11111: out = {   in[0],31'b0};
			
			// Shift Right Logical
			7'b01_00000: out = in[31:0];
			7'b01_00001: out = {1'b0, in[31:1] };
			7'b01_00010: out = {2'b0, in[31:2] };
			7'b01_00011: out = {3'b0, in[31:3] };
			7'b01_00100: out = {4'b0, in[31:4] };
			7'b01_00101: out = {5'b0, in[31:5] };
			7'b01_00110: out = {6'b0, in[31:6] };
			7'b01_00111: out = {7'b0, in[31:7] };
			7'b01_01000: out = {8'b0, in[31:8] };
			7'b01_01001: out = {9'b0, in[31:9] };
			7'b01_01010: out = {10'b0,in[31:10]};
			7'b01_01011: out = {11'b0,in[31:11]};
			7'b01_01100: out = {12'b0,in[31:12]};
			7'b01_01101: out = {13'b0,in[31:13]};
			7'b01_01110: out = {14'b0,in[31:14]};
			7'b01_01111: out = {15'b0,in[31:15]};
			7'b01_10000: out = {16'b0,in[31:16]};
			7'b01_10001: out = {17'b0,in[31:17]};
			7'b01_10010: out = {18'b0,in[31:18]};
			7'b01_10011: out = {19'b0,in[31:19]};
			7'b01_10100: out = {20'b0,in[31:20]};
			7'b01_10101: out = {21'b0,in[31:21]};
			7'b01_10110: out = {22'b0,in[31:22]};
			7'b01_10111: out = {23'b0,in[31:23]};
			7'b01_11000: out = {24'b0,in[31:24]};
			7'b01_11001: out = {25'b0,in[31:25]};
			7'b01_11010: out = {26'b0,in[31:26]};
			7'b01_11011: out = {27'b0,in[31:27]};
			7'b01_11100: out = {28'b0,in[31:28]};
			7'b01_11101: out = {29'b0,in[31:29]};
			7'b01_11110: out = {30'b0,in[31:30]};
			7'b01_11111: out = {31'b0,in[31]};
			
			// Shift Right Arithmetic
			7'b10_00000: out = in[31:0];
			7'b10_00001: out = {in[31],in[31:1]       };
			7'b10_00010: out = {{2{in[31]}} ,in[31:2] };
			7'b10_00011: out = {{3{in[31]}} ,in[31:3] };
			7'b10_00100: out = {{4{in[31]}} ,in[31:4] };
			7'b10_00101: out = {{5{in[31]}} ,in[31:5] };
			7'b10_00110: out = {{6{in[31]}} ,in[31:6] };
			7'b10_00111: out = {{7{in[31]}} ,in[31:7] };
			7'b10_01000: out = {{8{in[31]}} ,in[31:8] };
			7'b10_01001: out = {{9{in[31]}} ,in[31:9] };
			7'b10_01010: out = {{10{in[31]}},in[31:10]};
			7'b10_01011: out = {{11{in[31]}},in[31:11]};
			7'b10_01100: out = {{12{in[31]}},in[31:12]};
			7'b10_01101: out = {{13{in[31]}},in[31:13]};
			7'b10_01110: out = {{14{in[31]}},in[31:14]};
			7'b10_01111: out = {{15{in[31]}},in[31:15]};
			7'b10_10000: out = {{16{in[31]}},in[31:16]};
			7'b10_10001: out = {{17{in[31]}},in[31:17]};
			7'b10_10010: out = {{18{in[31]}},in[31:18]};
			7'b10_10011: out = {{19{in[31]}},in[31:19]};
			7'b10_10100: out = {{20{in[31]}},in[31:20]};
			7'b10_10101: out = {{21{in[31]}},in[31:21]};
			7'b10_10110: out = {{22{in[31]}},in[31:22]};
			7'b10_10111: out = {{23{in[31]}},in[31:23]};
			7'b10_11000: out = {{24{in[31]}},in[31:24]};
			7'b10_11001: out = {{25{in[31]}},in[31:25]};
			7'b10_11010: out = {{26{in[31]}},in[31:26]};
			7'b10_11011: out = {{27{in[31]}},in[31:27]};
			7'b10_11100: out = {{28{in[31]}},in[31:28]};
			7'b10_11101: out = {{29{in[31]}},in[31:29]};
			7'b10_11110: out = {{30{in[31]}},in[31:30]};
			7'b10_11111: out = {{31{in[31]}},in[31]   };
			
			default: out = in;
		endcase
	end

endmodule
